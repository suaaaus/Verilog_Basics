module fa_v2 (a, b, ci, s);
input a, b, ci;
output s;

assign s=a^b^ci;


endmodule
